module hello(
	input clk);

initial
begin: proc_disp_hi
	$display("Hello");
end

endmodule
