package el2_lockstep_pkg;
  import el2_pkg::*;
  `include "el2_param.vh"
  ;//
  // Outputs
  typedef struct packed {
    logic                                 core_rst_l;
    logic [31:0]                          trace_rv_i_insn_ip;
    logic [31:0]                          trace_rv_i_address_ip;
    logic                                 trace_rv_i_valid_ip;
    logic                                 trace_rv_i_exception_ip;
    logic [4:0]                           trace_rv_i_ecause_ip;
    logic                                 trace_rv_i_interrupt_ip;
    logic [31:0]                          trace_rv_i_tval_ip;
    logic                                 dccm_clk_override;
    logic                                 icm_clk_override;
    logic                                 dec_tlu_core_ecc_disable;
    logic                                 o_cpu_halt_ack;
    logic                                 o_cpu_halt_status;
    logic                                 o_cpu_run_ack;
    logic                                 o_debug_mode_status;
    logic                                 mpc_debug_halt_ack;
    logic                                 mpc_debug_run_ack;
    logic                                 debug_brkpt_status;
    logic                                 dec_tlu_perfcnt0;
    logic                                 dec_tlu_perfcnt1;
    logic                                 dec_tlu_perfcnt2;
    logic                                 dec_tlu_perfcnt3;
    logic                                 dccm_wren;
    logic                                 dccm_rden;
    logic [pt.DCCM_BITS-1:0]              dccm_wr_addr_lo;
    logic [pt.DCCM_BITS-1:0]              dccm_wr_addr_hi;
    logic [pt.DCCM_BITS-1:0]              dccm_rd_addr_lo;
    logic [pt.DCCM_BITS-1:0]              dccm_rd_addr_hi;
    logic [pt.DCCM_FDATA_WIDTH-1:0]       dccm_wr_data_lo;
    logic [pt.DCCM_FDATA_WIDTH-1:0]       dccm_wr_data_hi;
    logic [pt.ICCM_BITS-1:1]              iccm_rw_addr;
    logic                                 iccm_wren;
    logic                                 iccm_rden;
    logic [2:0]                           iccm_wr_size;
    logic [77:0]                          iccm_wr_data;
    logic                                 iccm_buf_correct_ecc;
    logic                                 iccm_correction_state;
    logic [31:1]                          ic_rw_addr;
    logic [pt.ICACHE_NUM_WAYS-1:0]        ic_tag_valid;
    logic [pt.ICACHE_NUM_WAYS-1:0]        ic_wr_en;
    logic                                 ic_rd_en;
    logic [pt.ICACHE_BANKS_WAY-1:0][70:0] ic_wr_data;
    logic [70:0]                          ic_debug_wr_data;
    logic [63:0]                          ic_premux_data;
    logic                                 ic_sel_premux_data;
    logic [pt.ICACHE_INDEX_HI:3]          ic_debug_addr;
    logic                                 ic_debug_rd_en;
    logic                                 ic_debug_wr_en;
    logic                                 ic_debug_tag_array;
    logic [pt.ICACHE_NUM_WAYS-1:0]        ic_debug_way;
    logic                                 lsu_axi_awvalid;
    logic [pt.LSU_BUS_TAG-1:0]            lsu_axi_awid;
    logic [31:0]                          lsu_axi_awaddr;
    logic [3:0]                           lsu_axi_awregion;
    logic [7:0]                           lsu_axi_awlen;
    logic [2:0]                           lsu_axi_awsize;
    logic [1:0]                           lsu_axi_awburst;
    logic                                 lsu_axi_awlock;
    logic [3:0]                           lsu_axi_awcache;
    logic [2:0]                           lsu_axi_awprot;
    logic [3:0]                           lsu_axi_awqos;
    logic                                 lsu_axi_wvalid;
    logic [63:0]                          lsu_axi_wdata;
    logic [7:0]                           lsu_axi_wstrb;
    logic                                 lsu_axi_wlast;
    logic                                 lsu_axi_bready;
    logic                                 lsu_axi_arvalid;
    logic [pt.LSU_BUS_TAG-1:0]            lsu_axi_arid;
    logic [31:0]                          lsu_axi_araddr;
    logic [3:0]                           lsu_axi_arregion;
    logic [7:0]                           lsu_axi_arlen;
    logic [2:0]                           lsu_axi_arsize;
    logic [1:0]                           lsu_axi_arburst;
    logic                                 lsu_axi_arlock;
    logic [3:0]                           lsu_axi_arcache;
    logic [2:0]                           lsu_axi_arprot;
    logic [3:0]                           lsu_axi_arqos;
    logic                                 lsu_axi_rready;
    logic                                 ifu_axi_awvalid;
    logic [pt.IFU_BUS_TAG-1:0]            ifu_axi_awid;
    logic [31:0]                          ifu_axi_awaddr;
    logic [3:0]                           ifu_axi_awregion;
    logic [7:0]                           ifu_axi_awlen;
    logic [2:0]                           ifu_axi_awsize;
    logic [1:0]                           ifu_axi_awburst;
    logic                                 ifu_axi_awlock;
    logic [3:0]                           ifu_axi_awcache;
    logic [2:0]                           ifu_axi_awprot;
    logic [3:0]                           ifu_axi_awqos;
    logic                                 ifu_axi_wvalid;
    logic [63:0]                          ifu_axi_wdata;
    logic [7:0]                           ifu_axi_wstrb;
    logic                                 ifu_axi_wlast;
    logic                                 ifu_axi_bready;
    logic                                 ifu_axi_arvalid;
    logic [pt.IFU_BUS_TAG-1:0]            ifu_axi_arid;
    logic [31:0]                          ifu_axi_araddr;
    logic [3:0]                           ifu_axi_arregion;
    logic [7:0]                           ifu_axi_arlen;
    logic [2:0]                           ifu_axi_arsize;
    logic [1:0]                           ifu_axi_arburst;
    logic                                 ifu_axi_arlock;
    logic [3:0]                           ifu_axi_arcache;
    logic [2:0]                           ifu_axi_arprot;
    logic [3:0]                           ifu_axi_arqos;
    logic                                 ifu_axi_rready;
    logic                                 sb_axi_awvalid;
    logic [pt.SB_BUS_TAG-1:0]             sb_axi_awid;
    logic [31:0]                          sb_axi_awaddr;
    logic [3:0]                           sb_axi_awregion;
    logic [7:0]                           sb_axi_awlen;
    logic [2:0]                           sb_axi_awsize;
    logic [1:0]                           sb_axi_awburst;
    logic                                 sb_axi_awlock;
    logic [3:0]                           sb_axi_awcache;
    logic [2:0]                           sb_axi_awprot;
    logic [3:0]                           sb_axi_awqos;
    logic                                 sb_axi_wvalid;
    logic [63:0]                          sb_axi_wdata;
    logic [7:0]                           sb_axi_wstrb;
    logic                                 sb_axi_wlast;
    logic                                 sb_axi_bready;
    logic                                 sb_axi_arvalid;
    logic [pt.SB_BUS_TAG-1:0]             sb_axi_arid;
    logic [31:0]                          sb_axi_araddr;
    logic [3:0]                           sb_axi_arregion;
    logic [7:0]                           sb_axi_arlen;
    logic [2:0]                           sb_axi_arsize;
    logic [1:0]                           sb_axi_arburst;
    logic                                 sb_axi_arlock;
    logic [3:0]                           sb_axi_arcache;
    logic [2:0]                           sb_axi_arprot;
    logic [3:0]                           sb_axi_arqos;
    logic                                 sb_axi_rready;
    logic                                 dma_axi_awready;
    logic                                 dma_axi_wready;
    logic                                 dma_axi_bvalid;
    logic [1:0]                           dma_axi_bresp;
    logic [pt.DMA_BUS_TAG-1:0]            dma_axi_bid;
    logic                                 dma_axi_arready;
    logic                                 dma_axi_rvalid;
    logic [pt.DMA_BUS_TAG-1:0]            dma_axi_rid;
    logic [63:0]                          dma_axi_rdata;
    logic [1:0]                           dma_axi_rresp;
    logic                                 dma_axi_rlast;
    logic [31:0]                          haddr;
    logic [2:0]                           hburst;
    logic                                 hmastlock;
    logic [3:0]                           hprot;
    logic [2:0]                           hsize;
    logic [1:0]                           htrans;
    logic                                 hwrite;
    logic [31:0]                          lsu_haddr;
    logic [2:0]                           lsu_hburst;
    logic                                 lsu_hmastlock;
    logic [3:0]                           lsu_hprot;
    logic [2:0]                           lsu_hsize;
    logic [1:0]                           lsu_htrans;
    logic                                 lsu_hwrite;
    logic [63:0]                          lsu_hwdata;
    logic [31:0]                          sb_haddr;
    logic [2:0]                           sb_hburst;
    logic                                 sb_hmastlock;
    logic [3:0]                           sb_hprot;
    logic [2:0]                           sb_hsize;
    logic [1:0]                           sb_htrans;
    logic                                 sb_hwrite;
    logic [63:0]                          sb_hwdata;
    logic [63:0]                          dma_hrdata;
    logic                                 dma_hreadyout;
    logic                                 dma_hresp;
    logic [31:0]                          dmi_reg_rdata;
    logic                                 iccm_ecc_single_error;
    logic                                 iccm_ecc_double_error;
    logic                                 dccm_ecc_single_error;
    logic                                 dccm_ecc_double_error;
  } veer_outputs_t;

  // Inputs
  typedef struct packed {
    logic [31:1]                    rst_vec;
    logic                           nmi_int;
    logic [31:1]                    nmi_vec;
    logic                           i_cpu_halt_req;
    logic                           i_cpu_run_req;
    logic [31:4]                    core_id;
    logic                           mpc_debug_halt_req;
    logic                           mpc_debug_run_req;
    logic                           mpc_reset_run_req;
    logic [pt.DCCM_FDATA_WIDTH-1:0] dccm_rd_data_lo;
    logic [pt.DCCM_FDATA_WIDTH-1:0] dccm_rd_data_hi;
    logic [63:0]                    iccm_rd_data;
    logic [77:0]                    iccm_rd_data_ecc;
    logic [63:0]                    ic_rd_data;
    logic [70:0]                    ic_debug_rd_data;
    logic [25:0]                    ictag_debug_rd_data;
    logic [pt.ICACHE_BANKS_WAY-1:0] ic_eccerr;
    logic [pt.ICACHE_BANKS_WAY-1:0] ic_parerr;
    logic [pt.ICACHE_NUM_WAYS-1:0]  ic_rd_hit;
    logic                           ic_tag_perr;
    logic                           lsu_axi_awready;
    logic                           lsu_axi_wready;
    logic                           lsu_axi_bvalid;
    logic [1:0]                     lsu_axi_bresp;
    logic [pt.LSU_BUS_TAG-1:0]      lsu_axi_bid;
    logic                           lsu_axi_arready;
    logic                           lsu_axi_rvalid;
    logic [pt.LSU_BUS_TAG-1:0]      lsu_axi_rid;
    logic [63:0]                    lsu_axi_rdata;
    logic [1:0]                     lsu_axi_rresp;
    logic                           lsu_axi_rlast;
    logic                           ifu_axi_awready;
    logic                           ifu_axi_wready;
    logic                           ifu_axi_bvalid;
    logic [1:0]                     ifu_axi_bresp;
    logic [pt.IFU_BUS_TAG-1:0]      ifu_axi_bid;
    logic                           ifu_axi_arready;
    logic                           ifu_axi_rvalid;
    logic [pt.IFU_BUS_TAG-1:0]      ifu_axi_rid;
    logic [63:0]                    ifu_axi_rdata;
    logic [1:0]                     ifu_axi_rresp;
    logic                           ifu_axi_rlast;
    logic                           sb_axi_awready;
    logic                           sb_axi_wready;
    logic                           sb_axi_bvalid;
    logic [1:0]                     sb_axi_bresp;
    logic [pt.SB_BUS_TAG-1:0]       sb_axi_bid;
    logic                           sb_axi_arready;
    logic                           sb_axi_rvalid;
    logic [pt.SB_BUS_TAG-1:0]       sb_axi_rid;
    logic [63:0]                    sb_axi_rdata;
    logic [1:0]                     sb_axi_rresp;
    logic                           sb_axi_rlast;
    logic                           dma_axi_awvalid;
    logic [pt.DMA_BUS_TAG-1:0]      dma_axi_awid;
    logic [31:0]                    dma_axi_awaddr;
    logic [2:0]                     dma_axi_awsize;
    logic [2:0]                     dma_axi_awprot;
    logic [7:0]                     dma_axi_awlen;
    logic [1:0]                     dma_axi_awburst;
    logic                           dma_axi_wvalid;
    logic [63:0]                    dma_axi_wdata;
    logic [7:0]                     dma_axi_wstrb;
    logic                           dma_axi_wlast;
    logic                           dma_axi_bready;
    logic                           dma_axi_arvalid;
    logic [pt.DMA_BUS_TAG-1:0]      dma_axi_arid;
    logic [31:0]                    dma_axi_araddr;
    logic [2:0]                     dma_axi_arsize;
    logic [2:0]                     dma_axi_arprot;
    logic [7:0]                     dma_axi_arlen;
    logic [1:0]                     dma_axi_arburst;
    logic                           dma_axi_rready;
    logic [63:0]                    hrdata;
    logic                           hready;
    logic                           hresp;
    logic [63:0]                    lsu_hrdata;
    logic                           lsu_hready;
    logic                           lsu_hresp;
    logic [63:0]                    sb_hrdata;
    logic                           sb_hready;
    logic                           sb_hresp;
    logic                           dma_hsel;
    logic [31:0]                    dma_haddr;
    logic [2:0]                     dma_hburst;
    logic                           dma_hmastlock;
    logic [3:0]                     dma_hprot;
    logic [2:0]                     dma_hsize;
    logic [1:0]                     dma_htrans;
    logic                           dma_hwrite;
    logic [63:0]                    dma_hwdata;
    logic                           dma_hreadyin;
    logic                           lsu_bus_clk_en;
    logic                           ifu_bus_clk_en;
    logic                           dbg_bus_clk_en;
    logic                           dma_bus_clk_en;
    logic                           dmi_reg_en;
    logic [6:0]                     dmi_reg_addr;
    logic                           dmi_reg_wr_en;
    logic [31:0]                    dmi_reg_wdata;
    logic [pt.PIC_TOTAL_INT:1]      extintsrc_req;
    logic                           timer_int;
    logic                           soft_int;
    logic                           scan_mode;
  } veer_inputs_t;
endpackage
